`include "register_interface/typedef.svh"
`include "axi/typedef.svh"
`include "idma/typedef.svh"

/// iDMA top containing an AXI 64-bit descriptor based front-end and an AXI-Stream backend.
module idma_desc64fe_axisbe_wrap #(
    /// Width of the addresses
    parameter int unsigned AddrWidth              = 64   ,
    /// Width of a data item on the AXI bus
    parameter int unsigned DataWidth              = 64   ,
    /// Width an AXI ID
    parameter int unsigned AxiIdWidth             = 3    ,
    /// AXI user width
    parameter int unsigned UserWidth        = 32'd1,

    /// Specifies the depth of the fifo behind the descriptor address register
    parameter int unsigned InputFifoDepth   =     8,
    /// Specifies the buffer size of the fifo that tracks requests submitted to the backend
    parameter int unsigned PendingFifoDepth =     8,
    /// Specifies how many descriptors may be fetched speculatively
    parameter int unsigned NSpeculation     =     4,
     /// Number of transaction that can be in-flight concurrently
    parameter int unsigned NumAxInFlight    = 32'd3,
    /// The depth of the internal reorder buffer:
    /// - '2': minimal possible configuration
    /// - '3': efficiently handle misaligned transfers (recommended)
    parameter int unsigned BufferDepth      = 32'd2,
    /// How many requests the backend might have at the same time in its buffers.
    /// Usually, `NumAxInFlight + BufferDepth`
    parameter int unsigned BackendDepth     = NumAxInFlight + BufferDepth,
    /// With of a transfer: max transfer size is `2**TFLenWidth` bytes
    parameter int unsigned TFLenWidth       = 32'd32,
    /// The depth of the memory system the backend is attached to
    parameter int unsigned MemSysDepth      = 32'd0,
    /// Should both data shifts be done before the dataflow element?
    /// If this is enabled, then the data inserted into the dataflow element
    /// will no longer be word aligned, but only a single shifter is needed
    parameter bit          CombinedShifter  = 1'b0,
    /// Should the `R`-`AW` coupling hardware be present? (recommended)
    parameter bit          RAWCouplingAvail = 1'b0,
    /// Mask invalid data on the manager interface
    parameter bit MaskInvalidData            = 1'b1,
    /// Should hardware legalization be present? (recommended)
    /// If not, software legalization is required to ensure the transfers are
    /// AXI4-conformal
    parameter bit HardwareLegalizer          = 1'b1,
    /// Reject zero-length transfers
    parameter bit RejectZeroTransfers        = 1'b1,
    /// Should the error handler be present?
    parameter idma_pkg::error_cap_e ErrorCap = idma_pkg::NO_ERROR_HANDLING,
    /// Print the info of the FIFO configuration
    parameter bit PrintFifoInfo              = 1'b0,
    /// Strobe Width (do not override!)
    parameter int unsigned StrbWidth         = DataWidth / 8,
    /// Offset Width (do not override!)
    parameter int unsigned OffsetWidth       = $clog2(StrbWidth),
    /// AXI4+ATOP Request and Response channel type
    parameter type axi_req_t     = logic,
    parameter type axi_rsp_t     = logic,
    parameter type axi_r_chan_t  = logic,
    parameter type axi_w_chan_t  = logic,
    parameter type axi_ar_chan_t = logic,
    parameter type axi_aw_chan_t = logic,
    /// AXI Stream Request and Response channel type
    parameter type axis_req_t    = logic,
    parameter type axis_t_chan_t = logic,
    parameter type axis_rsp_t    = logic,
    /// regbus interface types. Use the REG_BUS_TYPEDEF macros to define the types
    /// or see the idma backend documentation for more details
    parameter type reg_rsp_t    = logic,
    parameter type reg_req_t    = logic
)(
    /// clock
    input  logic                  clk_i             ,
    /// reset
    input  logic                  rst_ni            ,
    /// Testmode in
    input  logic testmode_i,

    /// axi interface used for fetching descriptors from memory (frontend)
    /// master pair
    /// master request
    output axi_req_t              master_fe_req_o      ,
    /// master response
    input  axi_rsp_t              master_fe_rsp_i      ,
    /// ID to be used by the read channel
    input  logic [AxiIdWidth-1:0] axi_ar_id_i        ,
    /// ID to be used by the write channel
    input  logic [AxiIdWidth-1:0] axi_aw_id_i        ,
    /// AXI4 (slave) interface used for reg access.
    /// The slave interface exposes two registers: One address register to
    /// write a descriptor address to process and a status register that
    /// exposes whether the DMA is busy on bit 0 and whether FIFOs are full
    /// on bit 1.
    input  axi_req_t              slave_fe_req_i,
    output axi_rsp_t              slave_fe_rsp_o,

    // write axi stream interface used for backend connection
    output axis_req_t              streaming_wr_req_o,
    input  axis_rsp_t              streaming_wr_rsp_i,
    // read axi stream interface used for backend connection
    input  axis_req_t              streaming_rd_req_i,
    output axis_rsp_t              streaming_rd_rsp_o,

    // read/write axi master interface used for backend connection
    output axi_req_t master_be_axi_req_o,
    input  axi_rsp_t master_be_axi_rsp_i,

    /// Event: irq
    output logic                  irq_o
);

//-----------------------//
//  TYPE DEFINITIONS     //
//-----------------------//
localparam int unsigned OneDLength       = 32;
typedef logic [AddrWidth-1:0]  addr_t;
typedef logic [DataWidth-1:0]  data_t;
typedef logic [StrbWidth-1:0]  strb_t;
typedef logic [OneDLength-1:0] length_t;
typedef logic [AxiIdWidth-1:0] id_t;
typedef logic [UserWidth-1:0]  user_t;
typedef logic [TFLenWidth-1:0] tf_len_t;


typedef struct packed {
    axi_ar_chan_t ar_chan;
} axi_read_meta_channel_t;

typedef struct packed {
    axi_read_meta_channel_t axi;
} read_meta_channel_t;

typedef struct packed {
    axis_t_chan_t t_chan;
} axis_write_meta_channel_t;

typedef struct packed {
    axi_aw_chan_t aw_chan;
} axi_write_meta_channel_t;

typedef struct packed {
    axis_write_meta_channel_t axis;
    axi_write_meta_channel_t axi;
} write_meta_channel_t;

//--------------------------------------
// Connections between frontend and backend
//--------------------------------------
`IDMA_TYPEDEF_FULL_REQ_T(idma_req_t, id_t, addr_t, tf_len_t)
`IDMA_TYPEDEF_FULL_RSP_T(idma_rsp_t, addr_t)
// dma request
idma_req_t idma_req;
logic req_valid;
logic req_ready;

// dma response
idma_rsp_t idma_rsp;
logic rsp_valid;
logic rsp_ready;

// busy signal
idma_pkg::idma_busy_t busy;

///FRONT END AXI///
reg_req_t fe_reg_req;
reg_rsp_t fe_reg_rsp;

axi_to_reg_v2 #(
    .AxiAddrWidth   ( AddrWidth         ),
    .AxiDataWidth   ( DataWidth         ),
    .AxiIdWidth     ( AxiIdWidth        ),
    .AxiUserWidth   ( UserWidth         ),
    .RegDataWidth   ( DataWidth         ),
    .axi_req_t      ( axi_req_t         ),
    .axi_rsp_t      ( axi_rsp_t         ),
    .reg_req_t      ( reg_req_t         ),
    .reg_rsp_t      ( reg_rsp_t         )
) axi_to_reg (
    .clk_i          ( clk_i             ),
    .rst_ni         ( rst_ni            ),
    .axi_req_i      ( slave_fe_req_i    ),
    .axi_rsp_o      ( slave_fe_rsp_o    ),
    .reg_req_o      ( fe_reg_req        ),
    .reg_rsp_i      ( fe_reg_rsp        ),
    .reg_id_o       ( /*NOT USED*/      ),
    .busy_o         ( /*NOT USED*/      )
);

idma_desc64_top #(
    .AddrWidth        ( AddrWidth        ),
    .DataWidth        ( DataWidth        ),
    .AxiIdWidth       ( AxiIdWidth       ),
    .idma_req_t       ( idma_req_t       ),
    .idma_rsp_t       ( idma_rsp_t       ),
    .axi_req_t        ( axi_req_t        ),
    .axi_rsp_t        ( axi_rsp_t        ),
    .axi_ar_chan_t    ( axi_ar_chan_t    ),
    .axi_r_chan_t     ( axi_r_chan_t     ),
    .reg_req_t        ( reg_req_t        ),
    .reg_rsp_t        ( reg_rsp_t        ),
    .InputFifoDepth   ( InputFifoDepth   ),
    .PendingFifoDepth ( PendingFifoDepth ),
    .BackendDepth     ( BackendDepth ),
    .NSpeculation     ( NSpeculation )
) i_idma_frontend (
    .clk_i            ( clk_i           ),
    .rst_ni           ( rst_ni          ),
    .master_req_o     (master_fe_req_o ),
    .master_rsp_i     (master_fe_rsp_i ),
    .axi_ar_id_i      (axi_ar_id_i      ),
    .axi_aw_id_i      (axi_aw_id_i      ),
    .slave_req_i      (fe_reg_req       ),
    .slave_rsp_o      (fe_reg_rsp       ),
    .idma_req_o       (idma_req         ),
    .idma_req_valid_o (req_valid        ),
    .idma_req_ready_i (req_ready        ),
    .idma_rsp_i       (idma_rsp         ),
    .idma_rsp_valid_i (rsp_valid        ),
    .idma_rsp_ready_o (rsp_ready        ),
    .idma_busy_i      (|busy            ),
    .irq_o            (irq_o            )
);

axi_req_t be_axi_rd_req, be_axi_wr_req;
axi_rsp_t be_axi_rd_rsp, be_axi_wr_rsp;

///BACKEND AXI///
idma_backend_rw_axi_rw_axis #(
    .CombinedShifter      ( CombinedShifter      ),
    .DataWidth            ( DataWidth            ),
    .AddrWidth            ( AddrWidth            ),
    .AxiIdWidth           ( AxiIdWidth           ),
    .UserWidth            ( UserWidth            ),
    .TFLenWidth           ( TFLenWidth           ),
    .MaskInvalidData      ( MaskInvalidData      ),
    .BufferDepth          ( BufferDepth          ),
    .RAWCouplingAvail     ( RAWCouplingAvail     ),
    .HardwareLegalizer    ( HardwareLegalizer    ),
    .RejectZeroTransfers  ( RejectZeroTransfers  ),
    .ErrorCap             ( ErrorCap             ),
    .PrintFifoInfo        ( PrintFifoInfo        ),
    .NumAxInFlight        ( NumAxInFlight        ),
    .MemSysDepth          ( MemSysDepth          ),
    .idma_req_t           ( idma_req_t           ),
    .idma_rsp_t           ( idma_rsp_t           ),
    .idma_eh_req_t        ( idma_pkg::idma_eh_req_t),
    .idma_busy_t          ( idma_pkg::idma_busy_t),
    .axi_req_t ( axi_req_t ),
    .axi_rsp_t ( axi_rsp_t ),
    .axis_req_t ( axis_req_t ),
    .axis_rsp_t ( axis_rsp_t ),
    .write_meta_channel_t ( write_meta_channel_t ),
    .read_meta_channel_t  ( read_meta_channel_t  )
) i_idma_backend  (
    .clk_i                ( clk_i           ),
    .rst_ni               ( rst_ni          ),
    .testmode_i           ( testmode_i      ),
    .idma_req_i           ( idma_req        ),
    .req_valid_i          ( req_valid       ),
    .req_ready_o          ( req_ready       ),
    .idma_rsp_o           ( idma_rsp        ),
    .rsp_valid_o          ( rsp_valid       ),
    .rsp_ready_i          ( rsp_ready       ),
    .idma_eh_req_i        ( '0              ),
    .eh_req_valid_i       ( '0              ),
    .eh_req_ready_o       (                 ),
    .axi_read_req_o       ( be_axi_rd_req   ),
    .axi_read_rsp_i       ( be_axi_rd_rsp   ),
    .axis_read_req_i      (streaming_rd_req_i),
    .axis_read_rsp_o      (streaming_rd_rsp_o),
    .axi_write_req_o      ( be_axi_wr_req  ),
    .axi_write_rsp_i      ( be_axi_wr_rsp  ),
    .axis_write_req_o     (streaming_wr_req_o),
    .axis_write_rsp_i     (streaming_wr_rsp_i),
    .busy_o               ( busy            )
);

axi_rw_join #(
    .axi_req_t(axi_req_t),
    .axi_resp_t(axi_rsp_t)
) be_join (
    .clk_i              ( clk_i                 ),
    .rst_ni             ( rst_ni                ),
    
    .slv_read_req_i     ( be_axi_rd_req         ),
    .slv_read_resp_o     ( be_axi_rd_rsp         ),
    
    .slv_write_req_i    ( be_axi_wr_req         ),
    .slv_write_resp_o    ( be_axi_wr_rsp         ),
    
    .mst_req_o          ( master_be_axi_req_o   ),
    .mst_resp_i          ( master_be_axi_rsp_i   )
);

endmodule
